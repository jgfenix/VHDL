------- inicio do componente mux 2x1 ----------
library ieee;
use ieee.std_logic_1164.all;

entity mux2x1 is
	port (A: in bit; B: in bit; C: in bit; S: out bit);
end mux2x1;
------- fim do componente mux 2x1 ----------